module XOR(input wire X0, input wire X1, output wire Y);
    assign Y = X0 ^ X1;
endmodule
